library verilog;
use verilog.vl_types.all;
entity waiting_time_t is
end waiting_time_t;
