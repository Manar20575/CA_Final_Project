library verilog;
use verilog.vl_types.all;
entity unit_t is
end unit_t;
