library verilog;
use verilog.vl_types.all;
entity Teller_t is
end Teller_t;
