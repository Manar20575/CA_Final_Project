library verilog;
use verilog.vl_types.all;
entity flags_t is
end flags_t;
