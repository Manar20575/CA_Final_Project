library verilog;
use verilog.vl_types.all;
entity unit_test_t is
end unit_test_t;
