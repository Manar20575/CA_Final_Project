library verilog;
use verilog.vl_types.all;
entity seg_t is
end seg_t;
