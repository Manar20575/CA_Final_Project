library verilog;
use verilog.vl_types.all;
entity counter_t is
end counter_t;
