library verilog;
use verilog.vl_types.all;
entity teller_t is
end teller_t;
