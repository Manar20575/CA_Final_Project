library verilog;
use verilog.vl_types.all;
entity wtime_t is
end wtime_t;
